`timescale 1ns / 1ns

// 串口接收缓冲
module uart_fifo_rx(

    );
endmodule
