`timescale 1ns / 1ns

// 串口发送缓冲
module uart_fifo_tx(

    );
endmodule
