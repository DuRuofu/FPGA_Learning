`timescale 1ns / 1ns

// 按照 I2C 协议对 EERPROM 存储芯片执行数据读写操作

module i2c_ctrl(

    );
endmodule
